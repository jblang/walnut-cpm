Date: Wednesday, 26 June 1985
From: John Blalock
Re:   Anti-APS Circuit

Summertime and the summer showers and power outages are almost here again.
Most of us use the standard surge and/or transient suppressors to protect
our systems from power line problems, but I also recommend use of the
following circuit:


				ANTI-APS CIRCUIT


                                                                   AC HIGH
              / Main Switch                        ----------O------------->  
       ,----o/ o-----------------------o-----------/\            TO SYSTEM
       o       S1                      |                                   
      (_  Main                         |           ----------O-,           
  F1    ) Fuse                ,--------o-----------/\          |           
       o                      |            ,-------------------'           
       |          Momentary |_o S2         |      -------                  
To 120 |          Start     | o            o------|     | 120 VAC DPST-NO  
VAC    |          Switch      |            |      | K1  | RELAY            
  _  HI|                      '------------'      |     |----.             
-| \---'                                          -------    |             
=|  |---|> Chassis Ground                                    |     AC NEUT   
-|_/---------------------------------------------------------o------------->  
     NEUT                                                        TO SYSTEM

Closing S1 does not turn on AC to the system, it just enables the
circuit.  Once S1 is closed, closing momentary switch S2 energizes K1.
One set of contacts on K1 provides AC to the system, the other
contacts are in parallel with S2 and latch K1 on until S1 is opened or
the main AC source goes off momentarily.  You need this circuit if you
have a "public utility" known to have frequent, unpredictable, power
outages.  If there is a momentary power failure, your system will shut
down until you restart it by pressing S2.  This prevents frequent
up/down AC surges like we see in Phoenix from being seen by your
system.  Make sure that the current ratings of F1, S1, and K1 exceed
your requirements.

John Blalock, W7AAY

uucp:	 ...{amd,decvax,hao,ihnp4,seismo}!noao!terak!jb
phone:	 (602) 998-4800
us mail: Terak Corp., 14151 N. 76th St., Scottsdale, AZ 85260
         \\\\\
          -----> Soon to be part of CalComp, A Sanders Company
